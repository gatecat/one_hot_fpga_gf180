VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO N_term_single
  CLASS BLOCK ;
  FOREIGN N_term_single ;
  ORIGIN 0.000 0.000 ;
  SIZE 390.000 BY 180.000 ;
  PIN Ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 142.520 0.000 143.080 2.000 ;
    END
  END Ci
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 291.480 0.000 292.040 2.000 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 318.360 0.000 318.920 2.000 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 321.720 0.000 322.280 2.000 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 323.960 0.000 324.520 2.000 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 327.320 0.000 327.880 2.000 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.560 0.000 330.120 2.000 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 332.920 0.000 333.480 2.000 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 335.160 0.000 335.720 2.000 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 337.400 0.000 337.960 2.000 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 340.760 0.000 341.320 2.000 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 343.000 0.000 343.560 2.000 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 294.840 0.000 295.400 2.000 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 346.360 0.000 346.920 2.000 ;
    END
  END FrameStrobe[20]
  PIN FrameStrobe[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 348.600 0.000 349.160 2.000 ;
    END
  END FrameStrobe[21]
  PIN FrameStrobe[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 351.960 0.000 352.520 2.000 ;
    END
  END FrameStrobe[22]
  PIN FrameStrobe[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 354.200 0.000 354.760 2.000 ;
    END
  END FrameStrobe[23]
  PIN FrameStrobe[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 356.440 0.000 357.000 2.000 ;
    END
  END FrameStrobe[24]
  PIN FrameStrobe[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 359.800 0.000 360.360 2.000 ;
    END
  END FrameStrobe[25]
  PIN FrameStrobe[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 362.040 0.000 362.600 2.000 ;
    END
  END FrameStrobe[26]
  PIN FrameStrobe[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 365.400 0.000 365.960 2.000 ;
    END
  END FrameStrobe[27]
  PIN FrameStrobe[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 367.640 0.000 368.200 2.000 ;
    END
  END FrameStrobe[28]
  PIN FrameStrobe[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 371.000 0.000 371.560 2.000 ;
    END
  END FrameStrobe[29]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 297.080 0.000 297.640 2.000 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 373.240 0.000 373.800 2.000 ;
    END
  END FrameStrobe[30]
  PIN FrameStrobe[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 375.480 0.000 376.040 2.000 ;
    END
  END FrameStrobe[31]
  PIN FrameStrobe[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 378.840 0.000 379.400 2.000 ;
    END
  END FrameStrobe[32]
  PIN FrameStrobe[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 381.080 0.000 381.640 2.000 ;
    END
  END FrameStrobe[33]
  PIN FrameStrobe[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 384.440 0.000 385.000 2.000 ;
    END
  END FrameStrobe[34]
  PIN FrameStrobe[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 386.680 0.000 387.240 2.000 ;
    END
  END FrameStrobe[35]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 299.320 0.000 299.880 2.000 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 302.680 0.000 303.240 2.000 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 304.920 0.000 305.480 2.000 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 308.280 0.000 308.840 2.000 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 310.520 0.000 311.080 2.000 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 313.880 0.000 314.440 2.000 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 316.120 0.000 316.680 2.000 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 21.560 178.000 22.120 180.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 123.480 178.000 124.040 180.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 133.560 178.000 134.120 180.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 143.640 178.000 144.200 180.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 153.720 178.000 154.280 180.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 164.920 178.000 165.480 180.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 175.000 178.000 175.560 180.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 185.080 178.000 185.640 180.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 195.160 178.000 195.720 180.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 205.240 178.000 205.800 180.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 215.320 178.000 215.880 180.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 31.640 178.000 32.200 180.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 225.400 178.000 225.960 180.000 ;
    END
  END FrameStrobe_O[20]
  PIN FrameStrobe_O[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 236.600 178.000 237.160 180.000 ;
    END
  END FrameStrobe_O[21]
  PIN FrameStrobe_O[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 246.680 178.000 247.240 180.000 ;
    END
  END FrameStrobe_O[22]
  PIN FrameStrobe_O[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 256.760 178.000 257.320 180.000 ;
    END
  END FrameStrobe_O[23]
  PIN FrameStrobe_O[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 266.840 178.000 267.400 180.000 ;
    END
  END FrameStrobe_O[24]
  PIN FrameStrobe_O[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 276.920 178.000 277.480 180.000 ;
    END
  END FrameStrobe_O[25]
  PIN FrameStrobe_O[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 287.000 178.000 287.560 180.000 ;
    END
  END FrameStrobe_O[26]
  PIN FrameStrobe_O[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 297.080 178.000 297.640 180.000 ;
    END
  END FrameStrobe_O[27]
  PIN FrameStrobe_O[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 307.160 178.000 307.720 180.000 ;
    END
  END FrameStrobe_O[28]
  PIN FrameStrobe_O[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 318.360 178.000 318.920 180.000 ;
    END
  END FrameStrobe_O[29]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 41.720 178.000 42.280 180.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 328.440 178.000 329.000 180.000 ;
    END
  END FrameStrobe_O[30]
  PIN FrameStrobe_O[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 338.520 178.000 339.080 180.000 ;
    END
  END FrameStrobe_O[31]
  PIN FrameStrobe_O[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 348.600 178.000 349.160 180.000 ;
    END
  END FrameStrobe_O[32]
  PIN FrameStrobe_O[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 358.680 178.000 359.240 180.000 ;
    END
  END FrameStrobe_O[33]
  PIN FrameStrobe_O[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 368.760 178.000 369.320 180.000 ;
    END
  END FrameStrobe_O[34]
  PIN FrameStrobe_O[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 378.840 178.000 379.400 180.000 ;
    END
  END FrameStrobe_O[35]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 51.800 178.000 52.360 180.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 61.880 178.000 62.440 180.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 71.960 178.000 72.520 180.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 83.160 178.000 83.720 180.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 93.240 178.000 93.800 180.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 103.320 178.000 103.880 180.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 113.400 178.000 113.960 180.000 ;
    END
  END FrameStrobe_O[9]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1.400 0.000 1.960 2.000 ;
    END
  END N1END[0]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.640 0.000 4.200 2.000 ;
    END
  END N1END[1]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 5.880 0.000 6.440 2.000 ;
    END
  END N1END[2]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 9.240 0.000 9.800 2.000 ;
    END
  END N1END[3]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.880 0.000 34.440 2.000 ;
    END
  END N2END[0]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 36.120 0.000 36.680 2.000 ;
    END
  END N2END[1]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 38.360 0.000 38.920 2.000 ;
    END
  END N2END[2]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 41.720 0.000 42.280 2.000 ;
    END
  END N2END[3]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.960 0.000 44.520 2.000 ;
    END
  END N2END[4]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.320 0.000 47.880 2.000 ;
    END
  END N2END[5]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 49.560 0.000 50.120 2.000 ;
    END
  END N2END[6]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 52.920 0.000 53.480 2.000 ;
    END
  END N2END[7]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 11.480 0.000 12.040 2.000 ;
    END
  END N2MID[0]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 14.840 0.000 15.400 2.000 ;
    END
  END N2MID[1]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 17.080 0.000 17.640 2.000 ;
    END
  END N2MID[2]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 19.320 0.000 19.880 2.000 ;
    END
  END N2MID[3]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 22.680 0.000 23.240 2.000 ;
    END
  END N2MID[4]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 24.920 0.000 25.480 2.000 ;
    END
  END N2MID[5]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 28.280 0.000 28.840 2.000 ;
    END
  END N2MID[6]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 30.520 0.000 31.080 2.000 ;
    END
  END N2MID[7]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 55.160 0.000 55.720 2.000 ;
    END
  END N4END[0]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 82.040 0.000 82.600 2.000 ;
    END
  END N4END[10]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 85.400 0.000 85.960 2.000 ;
    END
  END N4END[11]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 87.640 0.000 88.200 2.000 ;
    END
  END N4END[12]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 91.000 0.000 91.560 2.000 ;
    END
  END N4END[13]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 93.240 0.000 93.800 2.000 ;
    END
  END N4END[14]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 95.480 0.000 96.040 2.000 ;
    END
  END N4END[15]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 57.400 0.000 57.960 2.000 ;
    END
  END N4END[1]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 60.760 0.000 61.320 2.000 ;
    END
  END N4END[2]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.000 0.000 63.560 2.000 ;
    END
  END N4END[3]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 66.360 0.000 66.920 2.000 ;
    END
  END N4END[4]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 68.600 0.000 69.160 2.000 ;
    END
  END N4END[5]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 71.960 0.000 72.520 2.000 ;
    END
  END N4END[6]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 74.200 0.000 74.760 2.000 ;
    END
  END N4END[7]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 76.440 0.000 77.000 2.000 ;
    END
  END N4END[8]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 79.800 0.000 80.360 2.000 ;
    END
  END N4END[9]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 98.840 0.000 99.400 2.000 ;
    END
  END NN4END[0]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 125.720 0.000 126.280 2.000 ;
    END
  END NN4END[10]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 129.080 0.000 129.640 2.000 ;
    END
  END NN4END[11]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 131.320 0.000 131.880 2.000 ;
    END
  END NN4END[12]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 133.560 0.000 134.120 2.000 ;
    END
  END NN4END[13]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 136.920 0.000 137.480 2.000 ;
    END
  END NN4END[14]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 139.160 0.000 139.720 2.000 ;
    END
  END NN4END[15]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 101.080 0.000 101.640 2.000 ;
    END
  END NN4END[1]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 104.440 0.000 105.000 2.000 ;
    END
  END NN4END[2]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 106.680 0.000 107.240 2.000 ;
    END
  END NN4END[3]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 110.040 0.000 110.600 2.000 ;
    END
  END NN4END[4]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 112.280 0.000 112.840 2.000 ;
    END
  END NN4END[5]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 114.520 0.000 115.080 2.000 ;
    END
  END NN4END[6]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 117.880 0.000 118.440 2.000 ;
    END
  END NN4END[7]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 120.120 0.000 120.680 2.000 ;
    END
  END NN4END[8]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 123.480 0.000 124.040 2.000 ;
    END
  END NN4END[9]
  PIN OutputEnable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 289.240 0.000 289.800 2.000 ;
    END
  END OutputEnable
  PIN OutputEnable_O
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 11.480 178.000 12.040 180.000 ;
    END
  END OutputEnable_O
  PIN S1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.760 0.000 145.320 2.000 ;
    END
  END S1BEG[0]
  PIN S1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 148.120 0.000 148.680 2.000 ;
    END
  END S1BEG[1]
  PIN S1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 150.360 0.000 150.920 2.000 ;
    END
  END S1BEG[2]
  PIN S1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 152.600 0.000 153.160 2.000 ;
    END
  END S1BEG[3]
  PIN S2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 155.960 0.000 156.520 2.000 ;
    END
  END S2BEG[0]
  PIN S2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 158.200 0.000 158.760 2.000 ;
    END
  END S2BEG[1]
  PIN S2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 161.560 0.000 162.120 2.000 ;
    END
  END S2BEG[2]
  PIN S2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 163.800 0.000 164.360 2.000 ;
    END
  END S2BEG[3]
  PIN S2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 167.160 0.000 167.720 2.000 ;
    END
  END S2BEG[4]
  PIN S2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 169.400 0.000 169.960 2.000 ;
    END
  END S2BEG[5]
  PIN S2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 171.640 0.000 172.200 2.000 ;
    END
  END S2BEG[6]
  PIN S2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 175.000 0.000 175.560 2.000 ;
    END
  END S2BEG[7]
  PIN S2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 177.240 0.000 177.800 2.000 ;
    END
  END S2BEGb[0]
  PIN S2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 180.600 0.000 181.160 2.000 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 182.840 0.000 183.400 2.000 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 186.200 0.000 186.760 2.000 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 188.440 0.000 189.000 2.000 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 190.680 0.000 191.240 2.000 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.040 0.000 194.600 2.000 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 196.280 0.000 196.840 2.000 ;
    END
  END S2BEGb[7]
  PIN S4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 199.640 0.000 200.200 2.000 ;
    END
  END S4BEG[0]
  PIN S4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 226.520 0.000 227.080 2.000 ;
    END
  END S4BEG[10]
  PIN S4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 228.760 0.000 229.320 2.000 ;
    END
  END S4BEG[11]
  PIN S4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 232.120 0.000 232.680 2.000 ;
    END
  END S4BEG[12]
  PIN S4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 234.360 0.000 234.920 2.000 ;
    END
  END S4BEG[13]
  PIN S4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 237.720 0.000 238.280 2.000 ;
    END
  END S4BEG[14]
  PIN S4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 239.960 0.000 240.520 2.000 ;
    END
  END S4BEG[15]
  PIN S4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 201.880 0.000 202.440 2.000 ;
    END
  END S4BEG[1]
  PIN S4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.120 0.000 204.680 2.000 ;
    END
  END S4BEG[2]
  PIN S4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 207.480 0.000 208.040 2.000 ;
    END
  END S4BEG[3]
  PIN S4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 209.720 0.000 210.280 2.000 ;
    END
  END S4BEG[4]
  PIN S4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 213.080 0.000 213.640 2.000 ;
    END
  END S4BEG[5]
  PIN S4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 215.320 0.000 215.880 2.000 ;
    END
  END S4BEG[6]
  PIN S4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.680 0.000 219.240 2.000 ;
    END
  END S4BEG[7]
  PIN S4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 220.920 0.000 221.480 2.000 ;
    END
  END S4BEG[8]
  PIN S4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 223.160 0.000 223.720 2.000 ;
    END
  END S4BEG[9]
  PIN SS4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 242.200 0.000 242.760 2.000 ;
    END
  END SS4BEG[0]
  PIN SS4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 270.200 0.000 270.760 2.000 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 272.440 0.000 273.000 2.000 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 275.800 0.000 276.360 2.000 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 278.040 0.000 278.600 2.000 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 280.280 0.000 280.840 2.000 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 283.640 0.000 284.200 2.000 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 245.560 0.000 246.120 2.000 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 247.800 0.000 248.360 2.000 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 251.160 0.000 251.720 2.000 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 253.400 0.000 253.960 2.000 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 256.760 0.000 257.320 2.000 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 259.000 0.000 259.560 2.000 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 261.240 0.000 261.800 2.000 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 264.600 0.000 265.160 2.000 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 266.840 0.000 267.400 2.000 ;
    END
  END SS4BEG[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 285.880 0.000 286.440 2.000 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1.400 178.000 1.960 180.000 ;
    END
  END UserCLKo
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 52.960 7.540 54.560 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 147.040 7.540 148.640 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 241.120 7.540 242.720 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 335.200 7.540 336.800 168.860 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 100.000 7.540 101.600 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 194.080 7.540 195.680 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 288.160 7.540 289.760 168.860 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 382.240 7.540 383.840 168.860 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 7.540 383.840 168.860 ;
      LAYER Metal2 ;
        RECT 2.260 177.700 11.180 178.500 ;
        RECT 12.340 177.700 21.260 178.500 ;
        RECT 22.420 177.700 31.340 178.500 ;
        RECT 32.500 177.700 41.420 178.500 ;
        RECT 42.580 177.700 51.500 178.500 ;
        RECT 52.660 177.700 61.580 178.500 ;
        RECT 62.740 177.700 71.660 178.500 ;
        RECT 72.820 177.700 82.860 178.500 ;
        RECT 84.020 177.700 92.940 178.500 ;
        RECT 94.100 177.700 103.020 178.500 ;
        RECT 104.180 177.700 113.100 178.500 ;
        RECT 114.260 177.700 123.180 178.500 ;
        RECT 124.340 177.700 133.260 178.500 ;
        RECT 134.420 177.700 143.340 178.500 ;
        RECT 144.500 177.700 153.420 178.500 ;
        RECT 154.580 177.700 164.620 178.500 ;
        RECT 165.780 177.700 174.700 178.500 ;
        RECT 175.860 177.700 184.780 178.500 ;
        RECT 185.940 177.700 194.860 178.500 ;
        RECT 196.020 177.700 204.940 178.500 ;
        RECT 206.100 177.700 215.020 178.500 ;
        RECT 216.180 177.700 225.100 178.500 ;
        RECT 226.260 177.700 236.300 178.500 ;
        RECT 237.460 177.700 246.380 178.500 ;
        RECT 247.540 177.700 256.460 178.500 ;
        RECT 257.620 177.700 266.540 178.500 ;
        RECT 267.700 177.700 276.620 178.500 ;
        RECT 277.780 177.700 286.700 178.500 ;
        RECT 287.860 177.700 296.780 178.500 ;
        RECT 297.940 177.700 306.860 178.500 ;
        RECT 308.020 177.700 318.060 178.500 ;
        RECT 319.220 177.700 328.140 178.500 ;
        RECT 329.300 177.700 338.220 178.500 ;
        RECT 339.380 177.700 348.300 178.500 ;
        RECT 349.460 177.700 358.380 178.500 ;
        RECT 359.540 177.700 368.460 178.500 ;
        RECT 369.620 177.700 378.540 178.500 ;
        RECT 379.700 177.700 386.820 178.500 ;
        RECT 1.820 2.300 386.820 177.700 ;
        RECT 2.260 0.090 3.340 2.300 ;
        RECT 4.500 0.090 5.580 2.300 ;
        RECT 6.740 0.090 8.940 2.300 ;
        RECT 10.100 0.090 11.180 2.300 ;
        RECT 12.340 0.090 14.540 2.300 ;
        RECT 15.700 0.090 16.780 2.300 ;
        RECT 17.940 0.090 19.020 2.300 ;
        RECT 20.180 0.090 22.380 2.300 ;
        RECT 23.540 0.090 24.620 2.300 ;
        RECT 25.780 0.090 27.980 2.300 ;
        RECT 29.140 0.090 30.220 2.300 ;
        RECT 31.380 0.090 33.580 2.300 ;
        RECT 34.740 0.090 35.820 2.300 ;
        RECT 36.980 0.090 38.060 2.300 ;
        RECT 39.220 0.090 41.420 2.300 ;
        RECT 42.580 0.090 43.660 2.300 ;
        RECT 44.820 0.090 47.020 2.300 ;
        RECT 48.180 0.090 49.260 2.300 ;
        RECT 50.420 0.090 52.620 2.300 ;
        RECT 53.780 0.090 54.860 2.300 ;
        RECT 56.020 0.090 57.100 2.300 ;
        RECT 58.260 0.090 60.460 2.300 ;
        RECT 61.620 0.090 62.700 2.300 ;
        RECT 63.860 0.090 66.060 2.300 ;
        RECT 67.220 0.090 68.300 2.300 ;
        RECT 69.460 0.090 71.660 2.300 ;
        RECT 72.820 0.090 73.900 2.300 ;
        RECT 75.060 0.090 76.140 2.300 ;
        RECT 77.300 0.090 79.500 2.300 ;
        RECT 80.660 0.090 81.740 2.300 ;
        RECT 82.900 0.090 85.100 2.300 ;
        RECT 86.260 0.090 87.340 2.300 ;
        RECT 88.500 0.090 90.700 2.300 ;
        RECT 91.860 0.090 92.940 2.300 ;
        RECT 94.100 0.090 95.180 2.300 ;
        RECT 96.340 0.090 98.540 2.300 ;
        RECT 99.700 0.090 100.780 2.300 ;
        RECT 101.940 0.090 104.140 2.300 ;
        RECT 105.300 0.090 106.380 2.300 ;
        RECT 107.540 0.090 109.740 2.300 ;
        RECT 110.900 0.090 111.980 2.300 ;
        RECT 113.140 0.090 114.220 2.300 ;
        RECT 115.380 0.090 117.580 2.300 ;
        RECT 118.740 0.090 119.820 2.300 ;
        RECT 120.980 0.090 123.180 2.300 ;
        RECT 124.340 0.090 125.420 2.300 ;
        RECT 126.580 0.090 128.780 2.300 ;
        RECT 129.940 0.090 131.020 2.300 ;
        RECT 132.180 0.090 133.260 2.300 ;
        RECT 134.420 0.090 136.620 2.300 ;
        RECT 137.780 0.090 138.860 2.300 ;
        RECT 140.020 0.090 142.220 2.300 ;
        RECT 143.380 0.090 144.460 2.300 ;
        RECT 145.620 0.090 147.820 2.300 ;
        RECT 148.980 0.090 150.060 2.300 ;
        RECT 151.220 0.090 152.300 2.300 ;
        RECT 153.460 0.090 155.660 2.300 ;
        RECT 156.820 0.090 157.900 2.300 ;
        RECT 159.060 0.090 161.260 2.300 ;
        RECT 162.420 0.090 163.500 2.300 ;
        RECT 164.660 0.090 166.860 2.300 ;
        RECT 168.020 0.090 169.100 2.300 ;
        RECT 170.260 0.090 171.340 2.300 ;
        RECT 172.500 0.090 174.700 2.300 ;
        RECT 175.860 0.090 176.940 2.300 ;
        RECT 178.100 0.090 180.300 2.300 ;
        RECT 181.460 0.090 182.540 2.300 ;
        RECT 183.700 0.090 185.900 2.300 ;
        RECT 187.060 0.090 188.140 2.300 ;
        RECT 189.300 0.090 190.380 2.300 ;
        RECT 191.540 0.090 193.740 2.300 ;
        RECT 194.900 0.090 195.980 2.300 ;
        RECT 197.140 0.090 199.340 2.300 ;
        RECT 200.500 0.090 201.580 2.300 ;
        RECT 202.740 0.090 203.820 2.300 ;
        RECT 204.980 0.090 207.180 2.300 ;
        RECT 208.340 0.090 209.420 2.300 ;
        RECT 210.580 0.090 212.780 2.300 ;
        RECT 213.940 0.090 215.020 2.300 ;
        RECT 216.180 0.090 218.380 2.300 ;
        RECT 219.540 0.090 220.620 2.300 ;
        RECT 221.780 0.090 222.860 2.300 ;
        RECT 224.020 0.090 226.220 2.300 ;
        RECT 227.380 0.090 228.460 2.300 ;
        RECT 229.620 0.090 231.820 2.300 ;
        RECT 232.980 0.090 234.060 2.300 ;
        RECT 235.220 0.090 237.420 2.300 ;
        RECT 238.580 0.090 239.660 2.300 ;
        RECT 240.820 0.090 241.900 2.300 ;
        RECT 243.060 0.090 245.260 2.300 ;
        RECT 246.420 0.090 247.500 2.300 ;
        RECT 248.660 0.090 250.860 2.300 ;
        RECT 252.020 0.090 253.100 2.300 ;
        RECT 254.260 0.090 256.460 2.300 ;
        RECT 257.620 0.090 258.700 2.300 ;
        RECT 259.860 0.090 260.940 2.300 ;
        RECT 262.100 0.090 264.300 2.300 ;
        RECT 265.460 0.090 266.540 2.300 ;
        RECT 267.700 0.090 269.900 2.300 ;
        RECT 271.060 0.090 272.140 2.300 ;
        RECT 273.300 0.090 275.500 2.300 ;
        RECT 276.660 0.090 277.740 2.300 ;
        RECT 278.900 0.090 279.980 2.300 ;
        RECT 281.140 0.090 283.340 2.300 ;
        RECT 284.500 0.090 285.580 2.300 ;
        RECT 286.740 0.090 288.940 2.300 ;
        RECT 290.100 0.090 291.180 2.300 ;
        RECT 292.340 0.090 294.540 2.300 ;
        RECT 295.700 0.090 296.780 2.300 ;
        RECT 297.940 0.090 299.020 2.300 ;
        RECT 300.180 0.090 302.380 2.300 ;
        RECT 303.540 0.090 304.620 2.300 ;
        RECT 305.780 0.090 307.980 2.300 ;
        RECT 309.140 0.090 310.220 2.300 ;
        RECT 311.380 0.090 313.580 2.300 ;
        RECT 314.740 0.090 315.820 2.300 ;
        RECT 316.980 0.090 318.060 2.300 ;
        RECT 319.220 0.090 321.420 2.300 ;
        RECT 322.580 0.090 323.660 2.300 ;
        RECT 324.820 0.090 327.020 2.300 ;
        RECT 328.180 0.090 329.260 2.300 ;
        RECT 330.420 0.090 332.620 2.300 ;
        RECT 333.780 0.090 334.860 2.300 ;
        RECT 336.020 0.090 337.100 2.300 ;
        RECT 338.260 0.090 340.460 2.300 ;
        RECT 341.620 0.090 342.700 2.300 ;
        RECT 343.860 0.090 346.060 2.300 ;
        RECT 347.220 0.090 348.300 2.300 ;
        RECT 349.460 0.090 351.660 2.300 ;
        RECT 352.820 0.090 353.900 2.300 ;
        RECT 355.060 0.090 356.140 2.300 ;
        RECT 357.300 0.090 359.500 2.300 ;
        RECT 360.660 0.090 361.740 2.300 ;
        RECT 362.900 0.090 365.100 2.300 ;
        RECT 366.260 0.090 367.340 2.300 ;
        RECT 368.500 0.090 370.700 2.300 ;
        RECT 371.860 0.090 372.940 2.300 ;
        RECT 374.100 0.090 375.180 2.300 ;
        RECT 376.340 0.090 378.540 2.300 ;
        RECT 379.700 0.090 380.780 2.300 ;
        RECT 381.940 0.090 384.140 2.300 ;
        RECT 385.300 0.090 386.380 2.300 ;
      LAYER Metal3 ;
        RECT 1.770 0.140 386.870 169.540 ;
  END
END N_term_single
END LIBRARY

