VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO E_IO
  CLASS BLOCK ;
  FOREIGN E_IO ;
  ORIGIN 0.000 0.000 ;
  SIZE 110.000 BY 390.000 ;
  PIN A_I_top
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 1.400 110.000 1.960 ;
    END
  END A_I_top
  PIN A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 18.200 110.000 18.760 ;
    END
  END A_O_top
  PIN A_T_top
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 9.240 110.000 9.800 ;
    END
  END A_T_top
  PIN A_config_C_bit0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 51.800 110.000 52.360 ;
    END
  END A_config_C_bit0
  PIN A_config_C_bit1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 59.640 110.000 60.200 ;
    END
  END A_config_C_bit1
  PIN A_config_C_bit2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 68.600 110.000 69.160 ;
    END
  END A_config_C_bit2
  PIN A_config_C_bit3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 76.440 110.000 77.000 ;
    END
  END A_config_C_bit3
  PIN B_I_top
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 26.040 110.000 26.600 ;
    END
  END B_I_top
  PIN B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 42.840 110.000 43.400 ;
    END
  END B_O_top
  PIN B_T_top
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 35.000 110.000 35.560 ;
    END
  END B_T_top
  PIN B_config_C_bit0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 85.400 110.000 85.960 ;
    END
  END B_config_C_bit0
  PIN B_config_C_bit1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 93.240 110.000 93.800 ;
    END
  END B_config_C_bit1
  PIN B_config_C_bit2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 102.200 110.000 102.760 ;
    END
  END B_config_C_bit2
  PIN B_config_C_bit3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 111.160 110.000 111.720 ;
    END
  END B_config_C_bit3
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1.400 2.000 1.960 ;
    END
  END E1END[0]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3.640 2.000 4.200 ;
    END
  END E1END[1]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 7.000 2.000 7.560 ;
    END
  END E1END[2]
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 10.360 2.000 10.920 ;
    END
  END E1END[3]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 37.240 2.000 37.800 ;
    END
  END E2END[0]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 40.600 2.000 41.160 ;
    END
  END E2END[1]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 42.840 2.000 43.400 ;
    END
  END E2END[2]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 46.200 2.000 46.760 ;
    END
  END E2END[3]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 49.560 2.000 50.120 ;
    END
  END E2END[4]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 52.920 2.000 53.480 ;
    END
  END E2END[5]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 55.160 2.000 55.720 ;
    END
  END E2END[6]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 58.520 2.000 59.080 ;
    END
  END E2END[7]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 12.600 2.000 13.160 ;
    END
  END E2MID[0]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 15.960 2.000 16.520 ;
    END
  END E2MID[1]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 19.320 2.000 19.880 ;
    END
  END E2MID[2]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 21.560 2.000 22.120 ;
    END
  END E2MID[3]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 24.920 2.000 25.480 ;
    END
  END E2MID[4]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 28.280 2.000 28.840 ;
    END
  END E2MID[5]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 31.640 2.000 32.200 ;
    END
  END E2MID[6]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 33.880 2.000 34.440 ;
    END
  END E2MID[7]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 110.040 2.000 110.600 ;
    END
  END E6END[0]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 140.280 2.000 140.840 ;
    END
  END E6END[10]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 143.640 2.000 144.200 ;
    END
  END E6END[11]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 113.400 2.000 113.960 ;
    END
  END E6END[1]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 116.760 2.000 117.320 ;
    END
  END E6END[2]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 119.000 2.000 119.560 ;
    END
  END E6END[3]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 122.360 2.000 122.920 ;
    END
  END E6END[4]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 125.720 2.000 126.280 ;
    END
  END E6END[5]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.960 2.000 128.520 ;
    END
  END E6END[6]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 131.320 2.000 131.880 ;
    END
  END E6END[7]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.680 2.000 135.240 ;
    END
  END E6END[8]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 136.920 2.000 137.480 ;
    END
  END E6END[9]
  PIN EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 61.880 2.000 62.440 ;
    END
  END EE4END[0]
  PIN EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 92.120 2.000 92.680 ;
    END
  END EE4END[10]
  PIN EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 95.480 2.000 96.040 ;
    END
  END EE4END[11]
  PIN EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 97.720 2.000 98.280 ;
    END
  END EE4END[12]
  PIN EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 101.080 2.000 101.640 ;
    END
  END EE4END[13]
  PIN EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 104.440 2.000 105.000 ;
    END
  END EE4END[14]
  PIN EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 106.680 2.000 107.240 ;
    END
  END EE4END[15]
  PIN EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 64.120 2.000 64.680 ;
    END
  END EE4END[1]
  PIN EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 67.480 2.000 68.040 ;
    END
  END EE4END[2]
  PIN EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.840 2.000 71.400 ;
    END
  END EE4END[3]
  PIN EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 74.200 2.000 74.760 ;
    END
  END EE4END[4]
  PIN EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 76.440 2.000 77.000 ;
    END
  END EE4END[5]
  PIN EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 79.800 2.000 80.360 ;
    END
  END EE4END[6]
  PIN EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 83.160 2.000 83.720 ;
    END
  END EE4END[7]
  PIN EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 85.400 2.000 85.960 ;
    END
  END EE4END[8]
  PIN EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 88.760 2.000 89.320 ;
    END
  END EE4END[9]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 292.600 2.000 293.160 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 322.840 2.000 323.400 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 326.200 2.000 326.760 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 328.440 2.000 329.000 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 331.800 2.000 332.360 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 335.160 2.000 335.720 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 337.400 2.000 337.960 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 340.760 2.000 341.320 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 344.120 2.000 344.680 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 347.480 2.000 348.040 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 349.720 2.000 350.280 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 294.840 2.000 295.400 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 353.080 2.000 353.640 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 356.440 2.000 357.000 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 358.680 2.000 359.240 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 362.040 2.000 362.600 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 365.400 2.000 365.960 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 368.760 2.000 369.320 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 371.000 2.000 371.560 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 374.360 2.000 374.920 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 377.720 2.000 378.280 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 379.960 2.000 380.520 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 298.200 2.000 298.760 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 383.320 2.000 383.880 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 386.680 2.000 387.240 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 301.560 2.000 302.120 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 304.920 2.000 305.480 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 307.160 2.000 307.720 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 310.520 2.000 311.080 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 313.880 2.000 314.440 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 316.120 2.000 316.680 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 319.480 2.000 320.040 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 119.000 110.000 119.560 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 204.120 110.000 204.680 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 211.960 110.000 212.520 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 220.920 110.000 221.480 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 228.760 110.000 229.320 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 237.720 110.000 238.280 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 245.560 110.000 246.120 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 254.520 110.000 255.080 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 262.360 110.000 262.920 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 271.320 110.000 271.880 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 279.160 110.000 279.720 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 127.960 110.000 128.520 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 288.120 110.000 288.680 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 297.080 110.000 297.640 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 304.920 110.000 305.480 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 313.880 110.000 314.440 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 321.720 110.000 322.280 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 330.680 110.000 331.240 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 338.520 110.000 339.080 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 347.480 110.000 348.040 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 355.320 110.000 355.880 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 364.280 110.000 364.840 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 135.800 110.000 136.360 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 372.120 110.000 372.680 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 381.080 110.000 381.640 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 144.760 110.000 145.320 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 152.600 110.000 153.160 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 161.560 110.000 162.120 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 169.400 110.000 169.960 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 178.360 110.000 178.920 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 186.200 110.000 186.760 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 108.000 195.160 110.000 195.720 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 7.000 0.000 7.560 2.000 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 35.000 0.000 35.560 2.000 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 38.360 0.000 38.920 2.000 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.600 0.000 41.160 2.000 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.960 0.000 44.520 2.000 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 46.200 0.000 46.760 2.000 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 49.560 0.000 50.120 2.000 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 51.800 0.000 52.360 2.000 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 55.160 0.000 55.720 2.000 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 58.520 0.000 59.080 2.000 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 60.760 0.000 61.320 2.000 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 9.240 0.000 9.800 2.000 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 64.120 0.000 64.680 2.000 ;
    END
  END FrameStrobe[20]
  PIN FrameStrobe[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 66.360 0.000 66.920 2.000 ;
    END
  END FrameStrobe[21]
  PIN FrameStrobe[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 69.720 0.000 70.280 2.000 ;
    END
  END FrameStrobe[22]
  PIN FrameStrobe[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 71.960 0.000 72.520 2.000 ;
    END
  END FrameStrobe[23]
  PIN FrameStrobe[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 75.320 0.000 75.880 2.000 ;
    END
  END FrameStrobe[24]
  PIN FrameStrobe[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.560 0.000 78.120 2.000 ;
    END
  END FrameStrobe[25]
  PIN FrameStrobe[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.920 0.000 81.480 2.000 ;
    END
  END FrameStrobe[26]
  PIN FrameStrobe[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 84.280 0.000 84.840 2.000 ;
    END
  END FrameStrobe[27]
  PIN FrameStrobe[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 86.520 0.000 87.080 2.000 ;
    END
  END FrameStrobe[28]
  PIN FrameStrobe[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 89.880 0.000 90.440 2.000 ;
    END
  END FrameStrobe[29]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 12.600 0.000 13.160 2.000 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 92.120 0.000 92.680 2.000 ;
    END
  END FrameStrobe[30]
  PIN FrameStrobe[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 95.480 0.000 96.040 2.000 ;
    END
  END FrameStrobe[31]
  PIN FrameStrobe[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.720 0.000 98.280 2.000 ;
    END
  END FrameStrobe[32]
  PIN FrameStrobe[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 101.080 0.000 101.640 2.000 ;
    END
  END FrameStrobe[33]
  PIN FrameStrobe[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 103.320 0.000 103.880 2.000 ;
    END
  END FrameStrobe[34]
  PIN FrameStrobe[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 106.680 0.000 107.240 2.000 ;
    END
  END FrameStrobe[35]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 14.840 0.000 15.400 2.000 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 18.200 0.000 18.760 2.000 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 20.440 0.000 21.000 2.000 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 23.800 0.000 24.360 2.000 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.040 0.000 26.600 2.000 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 29.400 0.000 29.960 2.000 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 32.760 0.000 33.320 2.000 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 7.000 388.000 7.560 390.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 35.000 388.000 35.560 390.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 38.360 388.000 38.920 390.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.600 388.000 41.160 390.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.960 388.000 44.520 390.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 46.200 388.000 46.760 390.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 49.560 388.000 50.120 390.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 51.800 388.000 52.360 390.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 55.160 388.000 55.720 390.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 58.520 388.000 59.080 390.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 60.760 388.000 61.320 390.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 9.240 388.000 9.800 390.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 64.120 388.000 64.680 390.000 ;
    END
  END FrameStrobe_O[20]
  PIN FrameStrobe_O[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 66.360 388.000 66.920 390.000 ;
    END
  END FrameStrobe_O[21]
  PIN FrameStrobe_O[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 69.720 388.000 70.280 390.000 ;
    END
  END FrameStrobe_O[22]
  PIN FrameStrobe_O[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 71.960 388.000 72.520 390.000 ;
    END
  END FrameStrobe_O[23]
  PIN FrameStrobe_O[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 75.320 388.000 75.880 390.000 ;
    END
  END FrameStrobe_O[24]
  PIN FrameStrobe_O[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.560 388.000 78.120 390.000 ;
    END
  END FrameStrobe_O[25]
  PIN FrameStrobe_O[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.920 388.000 81.480 390.000 ;
    END
  END FrameStrobe_O[26]
  PIN FrameStrobe_O[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 84.280 388.000 84.840 390.000 ;
    END
  END FrameStrobe_O[27]
  PIN FrameStrobe_O[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 86.520 388.000 87.080 390.000 ;
    END
  END FrameStrobe_O[28]
  PIN FrameStrobe_O[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 89.880 388.000 90.440 390.000 ;
    END
  END FrameStrobe_O[29]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 12.600 388.000 13.160 390.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 92.120 388.000 92.680 390.000 ;
    END
  END FrameStrobe_O[30]
  PIN FrameStrobe_O[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 95.480 388.000 96.040 390.000 ;
    END
  END FrameStrobe_O[31]
  PIN FrameStrobe_O[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.720 388.000 98.280 390.000 ;
    END
  END FrameStrobe_O[32]
  PIN FrameStrobe_O[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 101.080 388.000 101.640 390.000 ;
    END
  END FrameStrobe_O[33]
  PIN FrameStrobe_O[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 103.320 388.000 103.880 390.000 ;
    END
  END FrameStrobe_O[34]
  PIN FrameStrobe_O[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 106.680 388.000 107.240 390.000 ;
    END
  END FrameStrobe_O[35]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 14.840 388.000 15.400 390.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 18.200 388.000 18.760 390.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 20.440 388.000 21.000 390.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 23.800 388.000 24.360 390.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.040 388.000 26.600 390.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 29.400 388.000 29.960 390.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 32.760 388.000 33.320 390.000 ;
    END
  END FrameStrobe_O[9]
  PIN OutputEnable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.640 0.000 4.200 2.000 ;
    END
  END OutputEnable
  PIN OutputEnable_O
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.640 388.000 4.200 390.000 ;
    END
  END OutputEnable_O
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1.400 0.000 1.960 2.000 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1.400 388.000 1.960 390.000 ;
    END
  END UserCLKo
  PIN W1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 147.000 2.000 147.560 ;
    END
  END W1BEG[0]
  PIN W1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 149.240 2.000 149.800 ;
    END
  END W1BEG[1]
  PIN W1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 152.600 2.000 153.160 ;
    END
  END W1BEG[2]
  PIN W1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 155.960 2.000 156.520 ;
    END
  END W1BEG[3]
  PIN W2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 158.200 2.000 158.760 ;
    END
  END W2BEG[0]
  PIN W2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 161.560 2.000 162.120 ;
    END
  END W2BEG[1]
  PIN W2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 164.920 2.000 165.480 ;
    END
  END W2BEG[2]
  PIN W2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 168.280 2.000 168.840 ;
    END
  END W2BEG[3]
  PIN W2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 170.520 2.000 171.080 ;
    END
  END W2BEG[4]
  PIN W2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 173.880 2.000 174.440 ;
    END
  END W2BEG[5]
  PIN W2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 177.240 2.000 177.800 ;
    END
  END W2BEG[6]
  PIN W2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 179.480 2.000 180.040 ;
    END
  END W2BEG[7]
  PIN W2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 182.840 2.000 183.400 ;
    END
  END W2BEGb[0]
  PIN W2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 186.200 2.000 186.760 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 189.560 2.000 190.120 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 191.800 2.000 192.360 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 195.160 2.000 195.720 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 198.520 2.000 199.080 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 200.760 2.000 201.320 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 204.120 2.000 204.680 ;
    END
  END W2BEGb[7]
  PIN W6BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 255.640 2.000 256.200 ;
    END
  END W6BEG[0]
  PIN W6BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 285.880 2.000 286.440 ;
    END
  END W6BEG[10]
  PIN W6BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 289.240 2.000 289.800 ;
    END
  END W6BEG[11]
  PIN W6BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 259.000 2.000 259.560 ;
    END
  END W6BEG[1]
  PIN W6BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 262.360 2.000 262.920 ;
    END
  END W6BEG[2]
  PIN W6BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 264.600 2.000 265.160 ;
    END
  END W6BEG[3]
  PIN W6BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 267.960 2.000 268.520 ;
    END
  END W6BEG[4]
  PIN W6BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 271.320 2.000 271.880 ;
    END
  END W6BEG[5]
  PIN W6BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 273.560 2.000 274.120 ;
    END
  END W6BEG[6]
  PIN W6BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 276.920 2.000 277.480 ;
    END
  END W6BEG[7]
  PIN W6BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 280.280 2.000 280.840 ;
    END
  END W6BEG[8]
  PIN W6BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 283.640 2.000 284.200 ;
    END
  END W6BEG[9]
  PIN WW4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 207.480 2.000 208.040 ;
    END
  END WW4BEG[0]
  PIN WW4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 237.720 2.000 238.280 ;
    END
  END WW4BEG[10]
  PIN WW4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 241.080 2.000 241.640 ;
    END
  END WW4BEG[11]
  PIN WW4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 243.320 2.000 243.880 ;
    END
  END WW4BEG[12]
  PIN WW4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 246.680 2.000 247.240 ;
    END
  END WW4BEG[13]
  PIN WW4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 250.040 2.000 250.600 ;
    END
  END WW4BEG[14]
  PIN WW4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 253.400 2.000 253.960 ;
    END
  END WW4BEG[15]
  PIN WW4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 210.840 2.000 211.400 ;
    END
  END WW4BEG[1]
  PIN WW4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 213.080 2.000 213.640 ;
    END
  END WW4BEG[2]
  PIN WW4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 216.440 2.000 217.000 ;
    END
  END WW4BEG[3]
  PIN WW4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 219.800 2.000 220.360 ;
    END
  END WW4BEG[4]
  PIN WW4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 222.040 2.000 222.600 ;
    END
  END WW4BEG[5]
  PIN WW4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 225.400 2.000 225.960 ;
    END
  END WW4BEG[6]
  PIN WW4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 228.760 2.000 229.320 ;
    END
  END WW4BEG[7]
  PIN WW4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 232.120 2.000 232.680 ;
    END
  END WW4BEG[8]
  PIN WW4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 234.360 2.000 234.920 ;
    END
  END WW4BEG[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 17.960 7.540 19.560 380.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 42.040 7.540 43.640 380.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 66.120 7.540 67.720 380.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 90.200 7.540 91.800 380.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 30.000 7.540 31.600 380.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 54.080 7.540 55.680 380.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 78.160 7.540 79.760 380.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 102.240 7.540 103.840 380.540 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 7.540 108.550 380.540 ;
      LAYER Metal2 ;
        RECT 0.140 387.700 1.100 388.500 ;
        RECT 2.260 387.700 3.340 388.500 ;
        RECT 4.500 387.700 6.700 388.500 ;
        RECT 7.860 387.700 8.940 388.500 ;
        RECT 10.100 387.700 12.300 388.500 ;
        RECT 13.460 387.700 14.540 388.500 ;
        RECT 15.700 387.700 17.900 388.500 ;
        RECT 19.060 387.700 20.140 388.500 ;
        RECT 21.300 387.700 23.500 388.500 ;
        RECT 24.660 387.700 25.740 388.500 ;
        RECT 26.900 387.700 29.100 388.500 ;
        RECT 30.260 387.700 32.460 388.500 ;
        RECT 33.620 387.700 34.700 388.500 ;
        RECT 35.860 387.700 38.060 388.500 ;
        RECT 39.220 387.700 40.300 388.500 ;
        RECT 41.460 387.700 43.660 388.500 ;
        RECT 44.820 387.700 45.900 388.500 ;
        RECT 47.060 387.700 49.260 388.500 ;
        RECT 50.420 387.700 51.500 388.500 ;
        RECT 52.660 387.700 54.860 388.500 ;
        RECT 56.020 387.700 58.220 388.500 ;
        RECT 59.380 387.700 60.460 388.500 ;
        RECT 61.620 387.700 63.820 388.500 ;
        RECT 64.980 387.700 66.060 388.500 ;
        RECT 67.220 387.700 69.420 388.500 ;
        RECT 70.580 387.700 71.660 388.500 ;
        RECT 72.820 387.700 75.020 388.500 ;
        RECT 76.180 387.700 77.260 388.500 ;
        RECT 78.420 387.700 80.620 388.500 ;
        RECT 81.780 387.700 83.980 388.500 ;
        RECT 85.140 387.700 86.220 388.500 ;
        RECT 87.380 387.700 89.580 388.500 ;
        RECT 90.740 387.700 91.820 388.500 ;
        RECT 92.980 387.700 95.180 388.500 ;
        RECT 96.340 387.700 97.420 388.500 ;
        RECT 98.580 387.700 100.780 388.500 ;
        RECT 101.940 387.700 103.020 388.500 ;
        RECT 104.180 387.700 106.380 388.500 ;
        RECT 107.540 387.700 109.620 388.500 ;
        RECT 0.140 2.300 109.620 387.700 ;
        RECT 0.140 0.090 1.100 2.300 ;
        RECT 2.260 0.090 3.340 2.300 ;
        RECT 4.500 0.090 6.700 2.300 ;
        RECT 7.860 0.090 8.940 2.300 ;
        RECT 10.100 0.090 12.300 2.300 ;
        RECT 13.460 0.090 14.540 2.300 ;
        RECT 15.700 0.090 17.900 2.300 ;
        RECT 19.060 0.090 20.140 2.300 ;
        RECT 21.300 0.090 23.500 2.300 ;
        RECT 24.660 0.090 25.740 2.300 ;
        RECT 26.900 0.090 29.100 2.300 ;
        RECT 30.260 0.090 32.460 2.300 ;
        RECT 33.620 0.090 34.700 2.300 ;
        RECT 35.860 0.090 38.060 2.300 ;
        RECT 39.220 0.090 40.300 2.300 ;
        RECT 41.460 0.090 43.660 2.300 ;
        RECT 44.820 0.090 45.900 2.300 ;
        RECT 47.060 0.090 49.260 2.300 ;
        RECT 50.420 0.090 51.500 2.300 ;
        RECT 52.660 0.090 54.860 2.300 ;
        RECT 56.020 0.090 58.220 2.300 ;
        RECT 59.380 0.090 60.460 2.300 ;
        RECT 61.620 0.090 63.820 2.300 ;
        RECT 64.980 0.090 66.060 2.300 ;
        RECT 67.220 0.090 69.420 2.300 ;
        RECT 70.580 0.090 71.660 2.300 ;
        RECT 72.820 0.090 75.020 2.300 ;
        RECT 76.180 0.090 77.260 2.300 ;
        RECT 78.420 0.090 80.620 2.300 ;
        RECT 81.780 0.090 83.980 2.300 ;
        RECT 85.140 0.090 86.220 2.300 ;
        RECT 87.380 0.090 89.580 2.300 ;
        RECT 90.740 0.090 91.820 2.300 ;
        RECT 92.980 0.090 95.180 2.300 ;
        RECT 96.340 0.090 97.420 2.300 ;
        RECT 98.580 0.090 100.780 2.300 ;
        RECT 101.940 0.090 103.020 2.300 ;
        RECT 104.180 0.090 106.380 2.300 ;
        RECT 107.540 0.090 109.620 2.300 ;
      LAYER Metal3 ;
        RECT 2.300 386.380 109.670 387.380 ;
        RECT 0.090 384.180 109.670 386.380 ;
        RECT 2.300 383.020 109.670 384.180 ;
        RECT 0.090 381.940 109.670 383.020 ;
        RECT 0.090 380.820 107.700 381.940 ;
        RECT 2.300 380.780 107.700 380.820 ;
        RECT 2.300 379.660 109.670 380.780 ;
        RECT 0.090 378.580 109.670 379.660 ;
        RECT 2.300 377.420 109.670 378.580 ;
        RECT 0.090 375.220 109.670 377.420 ;
        RECT 2.300 374.060 109.670 375.220 ;
        RECT 0.090 372.980 109.670 374.060 ;
        RECT 0.090 371.860 107.700 372.980 ;
        RECT 2.300 371.820 107.700 371.860 ;
        RECT 2.300 370.700 109.670 371.820 ;
        RECT 0.090 369.620 109.670 370.700 ;
        RECT 2.300 368.460 109.670 369.620 ;
        RECT 0.090 366.260 109.670 368.460 ;
        RECT 2.300 365.140 109.670 366.260 ;
        RECT 2.300 365.100 107.700 365.140 ;
        RECT 0.090 363.980 107.700 365.100 ;
        RECT 0.090 362.900 109.670 363.980 ;
        RECT 2.300 361.740 109.670 362.900 ;
        RECT 0.090 359.540 109.670 361.740 ;
        RECT 2.300 358.380 109.670 359.540 ;
        RECT 0.090 357.300 109.670 358.380 ;
        RECT 2.300 356.180 109.670 357.300 ;
        RECT 2.300 356.140 107.700 356.180 ;
        RECT 0.090 355.020 107.700 356.140 ;
        RECT 0.090 353.940 109.670 355.020 ;
        RECT 2.300 352.780 109.670 353.940 ;
        RECT 0.090 350.580 109.670 352.780 ;
        RECT 2.300 349.420 109.670 350.580 ;
        RECT 0.090 348.340 109.670 349.420 ;
        RECT 2.300 347.180 107.700 348.340 ;
        RECT 0.090 344.980 109.670 347.180 ;
        RECT 2.300 343.820 109.670 344.980 ;
        RECT 0.090 341.620 109.670 343.820 ;
        RECT 2.300 340.460 109.670 341.620 ;
        RECT 0.090 339.380 109.670 340.460 ;
        RECT 0.090 338.260 107.700 339.380 ;
        RECT 2.300 338.220 107.700 338.260 ;
        RECT 2.300 337.100 109.670 338.220 ;
        RECT 0.090 336.020 109.670 337.100 ;
        RECT 2.300 334.860 109.670 336.020 ;
        RECT 0.090 332.660 109.670 334.860 ;
        RECT 2.300 331.540 109.670 332.660 ;
        RECT 2.300 331.500 107.700 331.540 ;
        RECT 0.090 330.380 107.700 331.500 ;
        RECT 0.090 329.300 109.670 330.380 ;
        RECT 2.300 328.140 109.670 329.300 ;
        RECT 0.090 327.060 109.670 328.140 ;
        RECT 2.300 325.900 109.670 327.060 ;
        RECT 0.090 323.700 109.670 325.900 ;
        RECT 2.300 322.580 109.670 323.700 ;
        RECT 2.300 322.540 107.700 322.580 ;
        RECT 0.090 321.420 107.700 322.540 ;
        RECT 0.090 320.340 109.670 321.420 ;
        RECT 2.300 319.180 109.670 320.340 ;
        RECT 0.090 316.980 109.670 319.180 ;
        RECT 2.300 315.820 109.670 316.980 ;
        RECT 0.090 314.740 109.670 315.820 ;
        RECT 2.300 313.580 107.700 314.740 ;
        RECT 0.090 311.380 109.670 313.580 ;
        RECT 2.300 310.220 109.670 311.380 ;
        RECT 0.090 308.020 109.670 310.220 ;
        RECT 2.300 306.860 109.670 308.020 ;
        RECT 0.090 305.780 109.670 306.860 ;
        RECT 2.300 304.620 107.700 305.780 ;
        RECT 0.090 302.420 109.670 304.620 ;
        RECT 2.300 301.260 109.670 302.420 ;
        RECT 0.090 299.060 109.670 301.260 ;
        RECT 2.300 297.940 109.670 299.060 ;
        RECT 2.300 297.900 107.700 297.940 ;
        RECT 0.090 296.780 107.700 297.900 ;
        RECT 0.090 295.700 109.670 296.780 ;
        RECT 2.300 294.540 109.670 295.700 ;
        RECT 0.090 293.460 109.670 294.540 ;
        RECT 2.300 292.300 109.670 293.460 ;
        RECT 0.090 290.100 109.670 292.300 ;
        RECT 2.300 288.980 109.670 290.100 ;
        RECT 2.300 288.940 107.700 288.980 ;
        RECT 0.090 287.820 107.700 288.940 ;
        RECT 0.090 286.740 109.670 287.820 ;
        RECT 2.300 285.580 109.670 286.740 ;
        RECT 0.090 284.500 109.670 285.580 ;
        RECT 2.300 283.340 109.670 284.500 ;
        RECT 0.090 281.140 109.670 283.340 ;
        RECT 2.300 280.020 109.670 281.140 ;
        RECT 2.300 279.980 107.700 280.020 ;
        RECT 0.090 278.860 107.700 279.980 ;
        RECT 0.090 277.780 109.670 278.860 ;
        RECT 2.300 276.620 109.670 277.780 ;
        RECT 0.090 274.420 109.670 276.620 ;
        RECT 2.300 273.260 109.670 274.420 ;
        RECT 0.090 272.180 109.670 273.260 ;
        RECT 2.300 271.020 107.700 272.180 ;
        RECT 0.090 268.820 109.670 271.020 ;
        RECT 2.300 267.660 109.670 268.820 ;
        RECT 0.090 265.460 109.670 267.660 ;
        RECT 2.300 264.300 109.670 265.460 ;
        RECT 0.090 263.220 109.670 264.300 ;
        RECT 2.300 262.060 107.700 263.220 ;
        RECT 0.090 259.860 109.670 262.060 ;
        RECT 2.300 258.700 109.670 259.860 ;
        RECT 0.090 256.500 109.670 258.700 ;
        RECT 2.300 255.380 109.670 256.500 ;
        RECT 2.300 255.340 107.700 255.380 ;
        RECT 0.090 254.260 107.700 255.340 ;
        RECT 2.300 254.220 107.700 254.260 ;
        RECT 2.300 253.100 109.670 254.220 ;
        RECT 0.090 250.900 109.670 253.100 ;
        RECT 2.300 249.740 109.670 250.900 ;
        RECT 0.090 247.540 109.670 249.740 ;
        RECT 2.300 246.420 109.670 247.540 ;
        RECT 2.300 246.380 107.700 246.420 ;
        RECT 0.090 245.260 107.700 246.380 ;
        RECT 0.090 244.180 109.670 245.260 ;
        RECT 2.300 243.020 109.670 244.180 ;
        RECT 0.090 241.940 109.670 243.020 ;
        RECT 2.300 240.780 109.670 241.940 ;
        RECT 0.090 238.580 109.670 240.780 ;
        RECT 2.300 237.420 107.700 238.580 ;
        RECT 0.090 235.220 109.670 237.420 ;
        RECT 2.300 234.060 109.670 235.220 ;
        RECT 0.090 232.980 109.670 234.060 ;
        RECT 2.300 231.820 109.670 232.980 ;
        RECT 0.090 229.620 109.670 231.820 ;
        RECT 2.300 228.460 107.700 229.620 ;
        RECT 0.090 226.260 109.670 228.460 ;
        RECT 2.300 225.100 109.670 226.260 ;
        RECT 0.090 222.900 109.670 225.100 ;
        RECT 2.300 221.780 109.670 222.900 ;
        RECT 2.300 221.740 107.700 221.780 ;
        RECT 0.090 220.660 107.700 221.740 ;
        RECT 2.300 220.620 107.700 220.660 ;
        RECT 2.300 219.500 109.670 220.620 ;
        RECT 0.090 217.300 109.670 219.500 ;
        RECT 2.300 216.140 109.670 217.300 ;
        RECT 0.090 213.940 109.670 216.140 ;
        RECT 2.300 212.820 109.670 213.940 ;
        RECT 2.300 212.780 107.700 212.820 ;
        RECT 0.090 211.700 107.700 212.780 ;
        RECT 2.300 211.660 107.700 211.700 ;
        RECT 2.300 210.540 109.670 211.660 ;
        RECT 0.090 208.340 109.670 210.540 ;
        RECT 2.300 207.180 109.670 208.340 ;
        RECT 0.090 204.980 109.670 207.180 ;
        RECT 2.300 203.820 107.700 204.980 ;
        RECT 0.090 201.620 109.670 203.820 ;
        RECT 2.300 200.460 109.670 201.620 ;
        RECT 0.090 199.380 109.670 200.460 ;
        RECT 2.300 198.220 109.670 199.380 ;
        RECT 0.090 196.020 109.670 198.220 ;
        RECT 2.300 194.860 107.700 196.020 ;
        RECT 0.090 192.660 109.670 194.860 ;
        RECT 2.300 191.500 109.670 192.660 ;
        RECT 0.090 190.420 109.670 191.500 ;
        RECT 2.300 189.260 109.670 190.420 ;
        RECT 0.090 187.060 109.670 189.260 ;
        RECT 2.300 185.900 107.700 187.060 ;
        RECT 0.090 183.700 109.670 185.900 ;
        RECT 2.300 182.540 109.670 183.700 ;
        RECT 0.090 180.340 109.670 182.540 ;
        RECT 2.300 179.220 109.670 180.340 ;
        RECT 2.300 179.180 107.700 179.220 ;
        RECT 0.090 178.100 107.700 179.180 ;
        RECT 2.300 178.060 107.700 178.100 ;
        RECT 2.300 176.940 109.670 178.060 ;
        RECT 0.090 174.740 109.670 176.940 ;
        RECT 2.300 173.580 109.670 174.740 ;
        RECT 0.090 171.380 109.670 173.580 ;
        RECT 2.300 170.260 109.670 171.380 ;
        RECT 2.300 170.220 107.700 170.260 ;
        RECT 0.090 169.140 107.700 170.220 ;
        RECT 2.300 169.100 107.700 169.140 ;
        RECT 2.300 167.980 109.670 169.100 ;
        RECT 0.090 165.780 109.670 167.980 ;
        RECT 2.300 164.620 109.670 165.780 ;
        RECT 0.090 162.420 109.670 164.620 ;
        RECT 2.300 161.260 107.700 162.420 ;
        RECT 0.090 159.060 109.670 161.260 ;
        RECT 2.300 157.900 109.670 159.060 ;
        RECT 0.090 156.820 109.670 157.900 ;
        RECT 2.300 155.660 109.670 156.820 ;
        RECT 0.090 153.460 109.670 155.660 ;
        RECT 2.300 152.300 107.700 153.460 ;
        RECT 0.090 150.100 109.670 152.300 ;
        RECT 2.300 148.940 109.670 150.100 ;
        RECT 0.090 147.860 109.670 148.940 ;
        RECT 2.300 146.700 109.670 147.860 ;
        RECT 0.090 145.620 109.670 146.700 ;
        RECT 0.090 144.500 107.700 145.620 ;
        RECT 2.300 144.460 107.700 144.500 ;
        RECT 2.300 143.340 109.670 144.460 ;
        RECT 0.090 141.140 109.670 143.340 ;
        RECT 2.300 139.980 109.670 141.140 ;
        RECT 0.090 137.780 109.670 139.980 ;
        RECT 2.300 136.660 109.670 137.780 ;
        RECT 2.300 136.620 107.700 136.660 ;
        RECT 0.090 135.540 107.700 136.620 ;
        RECT 2.300 135.500 107.700 135.540 ;
        RECT 2.300 134.380 109.670 135.500 ;
        RECT 0.090 132.180 109.670 134.380 ;
        RECT 2.300 131.020 109.670 132.180 ;
        RECT 0.090 128.820 109.670 131.020 ;
        RECT 2.300 127.660 107.700 128.820 ;
        RECT 0.090 126.580 109.670 127.660 ;
        RECT 2.300 125.420 109.670 126.580 ;
        RECT 0.090 123.220 109.670 125.420 ;
        RECT 2.300 122.060 109.670 123.220 ;
        RECT 0.090 119.860 109.670 122.060 ;
        RECT 2.300 118.700 107.700 119.860 ;
        RECT 0.090 117.620 109.670 118.700 ;
        RECT 2.300 116.460 109.670 117.620 ;
        RECT 0.090 114.260 109.670 116.460 ;
        RECT 2.300 113.100 109.670 114.260 ;
        RECT 0.090 112.020 109.670 113.100 ;
        RECT 0.090 110.900 107.700 112.020 ;
        RECT 2.300 110.860 107.700 110.900 ;
        RECT 2.300 109.740 109.670 110.860 ;
        RECT 0.090 107.540 109.670 109.740 ;
        RECT 2.300 106.380 109.670 107.540 ;
        RECT 0.090 105.300 109.670 106.380 ;
        RECT 2.300 104.140 109.670 105.300 ;
        RECT 0.090 103.060 109.670 104.140 ;
        RECT 0.090 101.940 107.700 103.060 ;
        RECT 2.300 101.900 107.700 101.940 ;
        RECT 2.300 100.780 109.670 101.900 ;
        RECT 0.090 98.580 109.670 100.780 ;
        RECT 2.300 97.420 109.670 98.580 ;
        RECT 0.090 96.340 109.670 97.420 ;
        RECT 2.300 95.180 109.670 96.340 ;
        RECT 0.090 94.100 109.670 95.180 ;
        RECT 0.090 92.980 107.700 94.100 ;
        RECT 2.300 92.940 107.700 92.980 ;
        RECT 2.300 91.820 109.670 92.940 ;
        RECT 0.090 89.620 109.670 91.820 ;
        RECT 2.300 88.460 109.670 89.620 ;
        RECT 0.090 86.260 109.670 88.460 ;
        RECT 2.300 85.100 107.700 86.260 ;
        RECT 0.090 84.020 109.670 85.100 ;
        RECT 2.300 82.860 109.670 84.020 ;
        RECT 0.090 80.660 109.670 82.860 ;
        RECT 2.300 79.500 109.670 80.660 ;
        RECT 0.090 77.300 109.670 79.500 ;
        RECT 2.300 76.140 107.700 77.300 ;
        RECT 0.090 75.060 109.670 76.140 ;
        RECT 2.300 73.900 109.670 75.060 ;
        RECT 0.090 71.700 109.670 73.900 ;
        RECT 2.300 70.540 109.670 71.700 ;
        RECT 0.090 69.460 109.670 70.540 ;
        RECT 0.090 68.340 107.700 69.460 ;
        RECT 2.300 68.300 107.700 68.340 ;
        RECT 2.300 67.180 109.670 68.300 ;
        RECT 0.090 64.980 109.670 67.180 ;
        RECT 2.300 63.820 109.670 64.980 ;
        RECT 0.090 62.740 109.670 63.820 ;
        RECT 2.300 61.580 109.670 62.740 ;
        RECT 0.090 60.500 109.670 61.580 ;
        RECT 0.090 59.380 107.700 60.500 ;
        RECT 2.300 59.340 107.700 59.380 ;
        RECT 2.300 58.220 109.670 59.340 ;
        RECT 0.090 56.020 109.670 58.220 ;
        RECT 2.300 54.860 109.670 56.020 ;
        RECT 0.090 53.780 109.670 54.860 ;
        RECT 2.300 52.660 109.670 53.780 ;
        RECT 2.300 52.620 107.700 52.660 ;
        RECT 0.090 51.500 107.700 52.620 ;
        RECT 0.090 50.420 109.670 51.500 ;
        RECT 2.300 49.260 109.670 50.420 ;
        RECT 0.090 47.060 109.670 49.260 ;
        RECT 2.300 45.900 109.670 47.060 ;
        RECT 0.090 43.700 109.670 45.900 ;
        RECT 2.300 42.540 107.700 43.700 ;
        RECT 0.090 41.460 109.670 42.540 ;
        RECT 2.300 40.300 109.670 41.460 ;
        RECT 0.090 38.100 109.670 40.300 ;
        RECT 2.300 36.940 109.670 38.100 ;
        RECT 0.090 35.860 109.670 36.940 ;
        RECT 0.090 34.740 107.700 35.860 ;
        RECT 2.300 34.700 107.700 34.740 ;
        RECT 2.300 33.580 109.670 34.700 ;
        RECT 0.090 32.500 109.670 33.580 ;
        RECT 2.300 31.340 109.670 32.500 ;
        RECT 0.090 29.140 109.670 31.340 ;
        RECT 2.300 27.980 109.670 29.140 ;
        RECT 0.090 26.900 109.670 27.980 ;
        RECT 0.090 25.780 107.700 26.900 ;
        RECT 2.300 25.740 107.700 25.780 ;
        RECT 2.300 24.620 109.670 25.740 ;
        RECT 0.090 22.420 109.670 24.620 ;
        RECT 2.300 21.260 109.670 22.420 ;
        RECT 0.090 20.180 109.670 21.260 ;
        RECT 2.300 19.060 109.670 20.180 ;
        RECT 2.300 19.020 107.700 19.060 ;
        RECT 0.090 17.900 107.700 19.020 ;
        RECT 0.090 16.820 109.670 17.900 ;
        RECT 2.300 15.660 109.670 16.820 ;
        RECT 0.090 13.460 109.670 15.660 ;
        RECT 2.300 12.300 109.670 13.460 ;
        RECT 0.090 11.220 109.670 12.300 ;
        RECT 2.300 10.100 109.670 11.220 ;
        RECT 2.300 10.060 107.700 10.100 ;
        RECT 0.090 8.940 107.700 10.060 ;
        RECT 0.090 7.860 109.670 8.940 ;
        RECT 2.300 6.700 109.670 7.860 ;
        RECT 0.090 4.500 109.670 6.700 ;
        RECT 2.300 3.340 109.670 4.500 ;
        RECT 0.090 2.260 109.670 3.340 ;
        RECT 2.300 1.100 107.700 2.260 ;
        RECT 0.090 0.140 109.670 1.100 ;
      LAYER Metal4 ;
        RECT 0.140 380.840 109.060 385.750 ;
        RECT 0.140 7.240 17.660 380.840 ;
        RECT 19.860 7.240 29.700 380.840 ;
        RECT 31.900 7.240 41.740 380.840 ;
        RECT 43.940 7.240 53.780 380.840 ;
        RECT 55.980 7.240 65.820 380.840 ;
        RECT 68.020 7.240 77.860 380.840 ;
        RECT 80.060 7.240 89.900 380.840 ;
        RECT 92.100 7.240 101.940 380.840 ;
        RECT 104.140 7.240 109.060 380.840 ;
        RECT 0.140 2.330 109.060 7.240 ;
  END
END E_IO
END LIBRARY

